*nmos varying vto

.include /home/vlsilab/UG_students_2018/t14y_tsmc_025_level1.txt

m1 vdd in 0 0 RITSUBN1 l=1u w=0.5u

v_dd vdd 0 3.3
v_in in 0 3.3

.dc v_dd 0 3.3 0.1 v_in 0 3.3 1
.dc v_in 0 3.3 0.1 v_dd 0 3.3 1

.control

foreach lamda 0.010 0.031 0.1
altermod m1 LAMBDA = $lamda
run
end

.endc

.control

foreach iter 1 2 3 4 5 6 
setplot dc$iter
plot -v_dd#branch
end
.endc

.end