magic
tech scmos
timestamp 1522412051
<< nwell >>
rect 10 21 41 49
<< polysilicon >>
rect 16 33 18 35
rect 32 33 34 35
rect 16 11 18 26
rect 32 23 34 26
rect 16 7 17 11
rect 16 6 18 7
rect 32 6 34 19
rect 16 1 18 3
rect 32 1 34 3
<< ndiffusion >>
rect 14 3 16 6
rect 18 3 32 6
rect 34 3 35 6
<< pdiffusion >>
rect 15 30 16 33
rect 12 26 16 30
rect 18 30 32 33
rect 18 26 23 30
rect 27 26 32 30
rect 34 30 35 33
rect 34 26 38 30
<< metal1 >>
rect 10 48 41 49
rect 10 46 23 48
rect 11 34 15 46
rect 27 46 41 48
rect 35 34 39 46
rect 23 25 27 26
rect 10 22 27 25
rect 10 7 13 22
rect 36 -8 39 3
rect 10 -11 40 -8
<< ntransistor >>
rect 16 3 18 6
rect 32 3 34 6
<< ptransistor >>
rect 16 26 18 33
rect 32 26 34 33
<< polycontact >>
rect 32 19 36 23
rect 17 7 21 11
<< ndcontact >>
rect 10 3 14 7
rect 35 3 39 7
<< pdcontact >>
rect 11 30 15 34
rect 23 26 27 30
rect 35 30 39 34
<< nsubstratencontact >>
rect 23 44 27 48
<< labels >>
rlabel metal1 11 20 11 20 3 z
rlabel polycontact 34 21 34 21 1 b
rlabel polycontact 19 9 19 9 1 a
rlabel metal1 22 -9 22 -9 1 vss
rlabel metal1 18 48 18 48 5 vdd
<< end >>
