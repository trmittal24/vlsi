* SPICE3 file created from aoi.ext - technology: scmos
.include /home/barun/vlsi/t14y_tsmc_025_level3.txt
M1000 vdd a a_n27_8# vdd cmosp w=20u l=2u
+  ad=144p pd=56u as=520p ps=132u
M1001 a_n27_8# b vdd vdd cmosp w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 z c a_n27_8# vdd cmosp w=20u l=2u
+  ad=220p pd=62u as=0p ps=0u
M1003 a_n13_n16# a vss 0 cmosn w=10u l=2u
+  ad=70p pd=34u as=240p ps=88u
M1004 z b a_n13_n16# 0 cmosn w=10u l=2u
+  ad=140p pd=48u as=0p ps=0u
M1005 vss c z 0 cmosn w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 vss 0 9.7fF
C1 z 0 3.9fF
C2 c 0 4.9fF
C3 b 0 4.9fF
C4 a 0 4.9fF
C5 vdd 0 2.4fF

v_dd vdd 0 5 
v_ss vss 0 0 
v_a a 0 DC 1 PULSE(0 5 0ns 0ns 0ns 20ns 40ns )
v_b b 0 DC 1 PULSE(0 5 0ns 0ns 0ns 40ns 80ns )
v_c c 0 DC 1 PULSE(0 5 0ns 0ns 0ns 80ns 160ns )

.tran 0.01ns 200ns 

.control
run
setplot tran1
plot a b+5 c+10 z+15
.endc

.end