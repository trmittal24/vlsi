*Study of Cmos Gates 


.include /home/tarun/ngspice/t14y_tsmc_025_level3.txt


mpa vatob v_inb v_dd v_dd cmosp w=2u l=1u
mpb vnor v_ina vatob vatob cmosp w=2u l=1u
mna vnor v_ina 0 0 cmosn w=1u l=1u
mnb vnor v_inb 0 0 cmosn w=1u l=1u
c1 vnor 0 0.1f

vdd v_dd 0 5
vina v_ina 0 5
vinb v_inb 0 0
vina v_ina  0 pulse(0 5 2n 0.1n 0.1n 2n 5n) 
vinb v_inb  0 pulse(0 5 1n 0.1n 0.1n 2n 5n) 

.dc vina 0 5 0.01
.tran 0.01ns 5n
 
.control
        //0.44u 

foreach iter 0.44u   
alter mna w = $iter
alter mnb w = $iter
run
end
.endc

.control
foreach iter 1
*plot -v_dd#branch
setplot tran$iter
plot v_ina v_inb+5 vnor+10
//plot -v_dd#branch
meas tran vdmax1 MAX vnor from=0n to =0.9n
meas tran vdmin MIN vnor from=2.2n to =2.7n
meas tran vdmax2 MAX vnor from=4.3n to =4.9n

let rise1 = vdmin + 0.9*(vdmax1 - vdmin)
let rise2 = vdmin + 0.1*(vdmax1 - vdmin) 
let rise3 = vdmin + 0.9*(vdmax2 - vdmin)
meas tran tfall trig vnor val=rise1 fall=1 targ vnor val=rise2 fall=1
meas tran trise trig vnor val=rise2 rise=last targ vnor val=rise3 rise=last

let v1=0.5*v(v_dd)
meas tran t1 when v_inb=v1 cross=1
meas tran t2 when v_inb=v1 cross=2
meas tran i_int integ vdd#branch from=t1 to=t2
let power=(0-i_int*5)/(t2-t1)
print power

meas tran iavg AVG vdd#branch from=0n to =4n
let pow = iavg*5
print 'pow'

let v2 = (vdmax1 + vdmin)/2
meas tran tx when v_inb = v2 cross=1
meas tran ty when vnor = v2 cross=1

let tphl = ty - tx
print 'tphl'

meas tran tx1 when v_ina = v2 cross=2
meas tran ty1 when vnor = v2 cross=2

let tplh = ty1 - tx1
print 'tplh'

let tp = (tplh + tphl)/2
print 'tp'

end
.endc

.control

foreach iter 1 
setplot dc$iter
plot vnor

let der_v = deriv(vnor)
meas dc vil find v_ina when der_v = -1 fall=last
meas dc voh find vnor when v_ina=vil rise=last
meas dc vih find v_ina when der_v = -1 rise=last
meas dc vol find vnor when v_ina=vih rise=last

let nmh = voh - vih
let nml = vil - vol
print 'nmh'
print 'nml'
end
.endc

.end