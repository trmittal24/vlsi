*nmos load inverter

.include /home/vlsilab/UG_students_2018/t14y_tsmc_025_level3.txt

mdriver vd vg 0 0 cmosn w=1u l=1u
mload vdd vdd vd 0 cmosn w=1u l=1u

v_dd vdd 0 3
*vin vg 0 5

v_g vg 0 dc 1 pulse(0 3 1n 0.05n 0.05n 2n 4n) 

.tran 0.01ns 9n
*.dc v_g 0 5 0.1
*.measure tran vd_max MAX vd from=0n to =4n
*.measure tran vd_min MIN vd from=0n to =4n
*.measure tran id_avg AVG v_dd#branch from=0n to =4n 

.control
foreach wid 8u 10u 15u
foreach widm1 1u 2u 2.5u
alter mload w = 10*$wid
alter mdriver w = 95*$widm1
run
end
end


.endc



.control



foreach t 1 2 3 4 5 6 7 8 9 
setplot tran$t
*setplot dc$t
*plot vd  deriv(vd)
*setplot dc$t
plot vg vd v_dd#branch
*plot -v_dd#branch

let v1=0.5*vdd
meas tran t1 when vg=v1 cross=1
meas tran t2 when vg=v1 cross=2
meas tran i_int integ i(v_dd) from=t1 to=t2
let power=(0-i_int*vdd)/(t2-t1)
print 'power'


meas tran vd_max MAX v(vd) from=0n to =0.8n
meas tran vd_min MIN v(vd) from=1n to =1.2n 

let val1 = vd_min+0.1*(vd_max-vd_min)
let val2 = vd_min + 0.9*(vd_max - vd_min) 

meas tran trise TRIG v(vd) VAL=val1 RISE=1 TARG V(vd) VAL=val2  RISE=1 
meas tran tfall TRIG v(vd) VAL=val1 FALL=1 TARG V(vd) VAL=val2  FALL=1
end

.endc


.end