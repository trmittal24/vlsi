*nmos load

.include /home/tarun/ngspice/t14y_tsmc_025_level3.txt

mp vout vin vdd vdd cmosp l=1u w=1u
mn vout vin 0 0 cmosn l=1u w=1u

v_dd vdd 0 5
v_in vin 0 5

.dc v_in 0 5 0.1
.tran 0 4n
v_in vin 0 pulse(0 5 1n 0.1n 0.1n 2n 4n) 


.control

foreach iter 0.149u 0.147u 0.145u
alter mp l = $iter
run
end
.endc

.control
foreach iter 1 2 3 
*plot -v_dd#branch
setplot tran$iter
plot vin vout
plot -v_dd#branch
meas tran vdmax1 MAX vout from=0n to =0.8n
meas tran vdmin MIN vout from=1.5n to =2n
meas tran vdmax2 MAX vout from=3.2n to =3.5n

let rise1 = vdmin + 0.9*(vdmax1 - vdmin)
let rise2 = vdmin + 0.1*(vdmax1 - vdmin) 
let rise3 = vdmin + 0.9*(vdmax2 - vdmin)
meas tran tfall trig vout val=rise1 fall=1 targ vout val=rise2 fall=1
meas tran trise trig vout val=rise2 rise=last targ vout val=rise3 rise=last

let v1=0.5*vdd
meas tran t1 when vin=v1 cross=1
meas tran t2 when vin=v1 cross=2
meas tran i_int integ v_dd#branch from=t1 to=t2
let power=(0-i_int*5)/(t2-t1)
print power

meas tran iavg AVG v_dd#branch from=0n to =4n
let pow = iavg*5
print 'pow'

let v2 = (vdmax1 + vdmin)/2
meas tran tx when vin = v2 cross=1
meas tran ty when vout = v2 cross=1

let tphl = ty - tx
print 'tphl'



end
.endc

.control

foreach iter 1 2 3
setplot dc$iter
plot vout

let der_v = deriv(vout)
meas dc vil find vin when der_v = -1 fall=last
meas dc voh find vout when vin=vil rise=last
meas dc vol find vin when der_v = -1 rise=last
meas dc vol find vout when vin=vol rise=last

let nmh = voh - vol
let nml = vil - vol
print 'nmh'
print 'nml'
end
.endc

.end