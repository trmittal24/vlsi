magic
tech scmos
timestamp 1522411587
<< nwell >>
rect -15 33 69 60
<< polysilicon >>
rect -6 55 -4 59
rect 5 55 7 57
rect 28 48 30 57
rect 50 48 52 58
rect -6 19 -4 38
rect 5 31 7 38
rect 28 31 30 38
rect 50 31 52 38
rect -6 15 -5 19
rect -6 13 -4 15
rect 5 13 7 27
rect 28 13 30 27
rect 50 13 52 27
rect -6 1 -4 5
rect 5 2 7 5
rect 28 2 30 5
rect 50 3 52 5
<< ndiffusion >>
rect -9 9 -6 13
rect -13 5 -6 9
rect -4 9 5 13
rect -4 5 -2 9
rect 2 5 5 9
rect 7 10 15 13
rect 19 10 28 13
rect 7 5 28 10
rect 30 9 50 13
rect 30 5 39 9
rect 43 5 50 9
rect 52 11 62 13
rect 52 5 66 11
<< pdiffusion >>
rect -13 42 -6 55
rect -9 38 -6 42
rect -4 52 -1 55
rect 3 52 5 55
rect -4 38 5 52
rect 7 48 19 55
rect 7 38 28 48
rect 30 38 50 48
rect 52 42 67 48
rect 52 38 62 42
rect 66 38 67 42
<< metal1 >>
rect -15 58 69 60
rect -15 56 63 58
rect 67 56 69 58
rect -13 13 -10 38
rect 62 21 65 38
rect 16 19 65 21
rect -1 18 65 19
rect -1 15 19 18
rect 15 14 19 15
rect 62 15 65 18
rect -2 4 2 5
rect -15 3 2 4
rect 39 3 43 5
rect -15 0 66 3
<< ntransistor >>
rect -6 5 -4 13
rect 5 5 7 13
rect 28 5 30 13
rect 50 5 52 13
<< ptransistor >>
rect -6 38 -4 55
rect 5 38 7 55
rect 28 38 30 48
rect 50 38 52 48
<< polycontact >>
rect 5 27 9 31
rect 28 27 32 31
rect 50 27 54 31
rect -5 15 -1 19
<< ndcontact >>
rect -13 9 -9 13
rect -2 5 2 9
rect 15 10 19 14
rect 39 5 43 9
rect 62 11 66 15
<< pdcontact >>
rect -13 38 -9 42
rect -1 52 3 56
rect 62 38 66 42
<< nsubstratencontact >>
rect 63 54 67 58
<< labels >>
rlabel metal1 -11 24 -11 24 3 z
rlabel polycontact 7 29 7 29 1 a
rlabel polycontact 30 29 30 29 1 b
rlabel polycontact 52 29 52 29 1 c
rlabel metal1 42 59 42 59 5 vdd
rlabel metal1 45 1 45 1 1 vss
rlabel metal1 63 26 63 26 1 zn
<< end >>
