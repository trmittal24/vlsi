* SPICE3 file created from nor2.ext - technology: scmos

.include t14y_tsmc_025_level3.txt


M1000 a_16_26# a vdd vdd pfet w=17u l=2u
+ ad=243p pd=70u as=78p ps=46u 
M1001 z b a_16_26# vdd pfet w=10u l=2u
+ ad=58p pd=34u as=0p ps=0u 
M1002 z a vss 0 nfet w=8u l=2u
+ ad=144p pd=52u as=72p ps=52u 
M1003 vss b z 0 nfet w=8u l=2u
+ ad=0p pd=0u as=0p ps=0u 
C0 vdd b 2.6fF
C1 vss 0 4.7fF
C2 b 0 4.4fF
C3 a 0 4.4fF

v_dd vdd 0 5
v_ss vss 0 0
vina a  0 pulse(0 5 0n 0.1n 0.1n 10n 20n) 
vinb b  0 pulse(0 5 5n 0.1n 0.1n 10n 20n) 

//.dc vina 0 5 0.01
.tran 0.01ns 50n

.control 
run 
setplot tran1
plot  z a b
.endc

.end