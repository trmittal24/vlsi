magic
tech scmos
timestamp 1520939803
<< nwell >>
rect 0 24 50 53
<< polysilicon >>
rect 6 41 8 43
rect 21 41 23 43
rect 41 34 43 43
rect 6 20 8 24
rect 21 21 23 24
rect 6 16 7 20
rect 6 12 8 16
rect 21 12 23 17
rect 41 21 43 24
rect 41 12 43 17
rect 6 0 8 4
rect 21 2 23 4
rect 41 2 43 4
<< ndiffusion >>
rect 2 8 6 12
rect 5 4 6 8
rect 8 8 21 12
rect 8 4 16 8
rect 20 4 21 8
rect 23 8 30 12
rect 34 8 41 12
rect 23 4 41 8
rect 43 8 47 12
rect 43 4 44 8
<< pdiffusion >>
rect 2 28 6 41
rect 4 24 6 28
rect 8 36 15 41
rect 19 36 21 41
rect 8 24 21 36
rect 23 34 32 41
rect 23 24 41 34
rect 43 28 48 34
rect 43 24 46 28
<< metal1 >>
rect 15 52 48 53
rect 15 50 30 52
rect 15 41 19 50
rect 34 50 48 52
rect 1 8 4 24
rect 7 24 46 27
rect 7 20 10 24
rect 31 12 34 24
rect 16 3 20 4
rect 44 3 48 4
rect 16 0 48 3
<< ntransistor >>
rect 6 4 8 12
rect 21 4 23 12
rect 41 4 43 12
<< ptransistor >>
rect 6 24 8 41
rect 21 24 23 41
rect 41 24 43 34
<< polycontact >>
rect 7 16 11 20
rect 19 17 23 21
rect 41 17 45 21
<< ndcontact >>
rect 1 4 5 8
rect 16 4 20 8
rect 30 8 34 12
rect 44 4 48 8
<< pdcontact >>
rect 0 24 4 28
rect 15 36 19 41
rect 46 24 50 28
<< nsubstratencontact >>
rect 30 48 34 52
<< labels >>
rlabel metal1 29 2 29 2 1 vss
rlabel metal1 25 52 25 52 5 vdd
rlabel polycontact 21 19 21 19 1 a
rlabel polycontact 43 19 43 19 1 b
rlabel metal1 32 19 32 19 1 zn
rlabel metal1 3 17 3 17 3 z
<< end >>
