* SPICE3 file created from dl.ext - technology: scmos
.include t14y_tsmc_025_level3.txt

M1000 vdd c cn vdd pfet w=9u l=2u
+ ad=174p pd=78u as=62p ps=34u 
M1001 da cn d vdd pfet w=17u l=2u
+ ad=168p pd=86u as=93p ps=52u 
M1002 vdd da a_7_n14# vdd pfet w=9u l=2u
+ ad=0p pd=0u as=40p ps=28u 
M1003 z a_7_n14# vdd vdd pfet w=9u l=2u
+ ad=117p pd=44u as=0p ps=0u 
M1004 da c z vdd pfet w=9u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1005 vss c cn Gnd nfet w=5u l=2u
+ ad=114p pd=68u as=40p ps=28u 
M1006 da c d Gnd nfet w=13u l=2u
+ ad=115p pd=70u as=69p ps=44u 
M1007 vss da a_7_n14# Gnd nfet w=5u l=2u
+ ad=0p pd=0u as=116p ps=54u 
M1008 z a_7_n14# vss Gnd nfet w=5u l=2u
+ ad=69p pd=38u as=0p ps=0u 
M1009 da cn z Gnd nfet w=5u l=2u
+ ad=0p pd=0u as=0p ps=0u 
C0 vdd cn 8.4fF
C1 vss cn 3.0fF
C2 vdd c 23.3fF
C3 vdd da 7.1fF
C4 vdd a_7_n14# 10.4fF
C5 vss 0 16.0fF
C6 z 0 2.3fF
C7 a_7_n14# 0 5.7fF
C8 da 0 11.8fF
C9 cn 0 24.1fF
C10 c 0 15.4fF


vdd vdd 0 5
vss vss 0 0 
v_gg_c d 0 PULSE(0 5 0n 0.1n 0.1n 25n 50n)
v_gg_d c 0 PULSE(5 0 12n 0.1n 0.1n 50n 100n)


.control
 tran 0.01n 200n
 plot (c + 15) (cn + 10) (d + 5) z
 
.endc

.end0