* SPICE3 file created from nd3.ext - technology: scmos
.include t14y_tsmc_025_level3.txt

M1000 z a vdd vdd pfet w=7u l=2u
+ ad=189p pd=82u as=182p ps=80u 
M1001 vdd b z vdd pfet w=7u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1002 z c vdd vdd pfet w=7u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1003 a_n16_n33# a vss 0 nfet w=4u l=2u
+ ad=72p pd=44u as=32p ps=24u 
M1004 a_4_n33# b a_n16_n33# 0 nfet w=4u l=2u
+ ad=72p pd=44u as=0p ps=0u 
M1005 z c a_4_n33# 0 nfet w=4u l=2u
+ ad=36p pd=26u as=0p ps=0u 
C0 a vdd 3.3fF
C1 vdd b 3.3fF
C2 vdd vdd 12.7fF
C3 vdd c 3.3fF
C4 vdd z 5.9fF
C5 vss 0 13.2fF
C6 z 0 4.7fF
C7 c 0 7.1fF
C8 b 0 7.1fF
C9 a 0 7.1fF

v_dd vdd 0 5
v_ss vss 0 0 
v_gg_cp a 0 PULSE(0 5 0 0.1n 0.1n 15n 30n)
v_gg_d b 0 PULSE(0 5 0 0.1n 0.1n 30n 60n)
v_gg_d1 c 0 PULSE(0 5 0 0.1n 0.1n 60n 120n)

.control
 tran 0.01n 120n
setplot tran1
 plot (a + 15) (b + 10) (c + 5) (z)
 
.endc

.end