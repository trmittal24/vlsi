magic
tech scmos
timestamp 1521537788
<< nwell >>
rect -23 19 4 40
rect 26 19 48 40
rect 26 -40 42 -19
<< metal1 >>
rect -31 37 13 40
rect 30 37 42 40
rect -31 -37 -28 37
rect -15 18 -12 22
rect 25 17 27 21
rect 61 17 63 21
rect 10 12 12 16
rect 46 12 48 16
rect -23 1 4 3
rect 28 1 40 3
rect -23 -3 12 1
rect 28 0 42 1
rect 30 -3 42 0
rect 55 -1 67 3
rect 19 -16 22 -12
rect 55 -16 58 -12
rect 4 -21 6 -17
rect 29 -21 44 -17
rect -31 -40 12 -37
rect 26 -40 38 -37
<< metal2 >>
rect 0 26 51 29
rect 0 23 4 26
rect -28 -17 -25 18
rect -11 10 -8 18
rect 12 10 15 12
rect -11 7 15 10
rect 27 0 30 17
rect 48 16 51 26
rect 67 17 69 21
rect 35 7 38 13
rect 35 4 54 7
rect 15 -3 30 0
rect 15 -12 18 -3
rect 51 -12 54 4
rect 66 -16 69 17
rect -28 -20 0 -17
<< m2contact >>
rect -25 15 -21 19
rect -12 18 -8 22
rect 0 19 4 23
rect 27 17 31 21
rect 63 17 67 21
rect 12 12 16 16
rect 35 13 39 17
rect 48 12 52 16
rect 15 -16 19 -12
rect 51 -16 55 -12
rect 0 -21 4 -17
rect 65 -20 69 -16
use ../lab6/cmos_inverter  cmos_inverter_0
timestamp 1519723961
transform 1 0 -15 0 1 15
box -8 -13 4 25
use nd2  nd2_0
timestamp 1520932602
transform 1 0 -10 0 1 -2
box 10 2 41 42
use nd2  nd2_3
timestamp 1520932602
transform -1 0 41 0 -1 2
box 10 2 41 42
use nd2  nd2_1
timestamp 1520932602
transform 1 0 26 0 1 -2
box 10 2 41 42
use nd2  nd2_2
timestamp 1520932602
transform -1 0 77 0 -1 2
box 10 2 41 42
<< end >>
