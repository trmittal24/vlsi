magic
tech scmos
timestamp 1522412814
<< nwell >>
rect -27 8 24 38
<< polysilicon >>
rect -15 28 -13 30
rect -6 28 -4 30
rect 10 28 12 30
rect -15 5 -13 8
rect -6 1 -4 8
rect 10 7 12 8
rect -15 -6 -13 1
rect -6 -6 -4 -3
rect 10 -6 12 3
rect -15 -18 -13 -16
rect -6 -18 -4 -16
rect 10 -18 12 -16
<< ndiffusion >>
rect -27 -10 -15 -6
rect -23 -14 -15 -10
rect -27 -16 -15 -14
rect -13 -16 -6 -6
rect -4 -10 10 -6
rect -4 -14 2 -10
rect 6 -14 10 -10
rect -4 -16 10 -14
rect 12 -10 24 -6
rect 12 -14 20 -10
rect 12 -16 24 -14
<< pdiffusion >>
rect -27 18 -15 28
rect -27 14 -23 18
rect -19 14 -15 18
rect -27 8 -15 14
rect -13 25 -12 28
rect -8 25 -6 28
rect -13 8 -6 25
rect -4 18 10 28
rect -4 14 -1 18
rect 3 14 10 18
rect -4 8 10 14
rect 12 18 23 28
rect 12 14 17 18
rect 21 14 23 18
rect 12 8 23 14
<< metal1 >>
rect -27 36 24 38
rect -27 33 2 36
rect -11 29 -8 33
rect 6 33 24 36
rect -19 14 -1 16
rect -22 13 2 14
rect 18 -1 21 14
rect 2 -4 21 -1
rect 2 -10 5 -4
rect -27 -17 -23 -14
rect 20 -17 24 -14
rect -27 -22 24 -17
<< ntransistor >>
rect -15 -16 -13 -6
rect -6 -16 -4 -6
rect 10 -16 12 -6
<< ptransistor >>
rect -15 8 -13 28
rect -6 8 -4 28
rect 10 8 12 28
<< polycontact >>
rect -16 1 -12 5
rect 10 3 14 7
rect -7 -3 -3 1
<< ndcontact >>
rect -27 -14 -23 -10
rect 2 -14 6 -10
rect 20 -14 24 -10
<< pdcontact >>
rect -23 14 -19 18
rect -12 25 -8 29
rect -1 14 3 18
rect 17 14 21 18
<< nsubstratencontact >>
rect 2 32 6 36
<< labels >>
rlabel polycontact -5 -1 -5 -1 1 b
rlabel polycontact 12 5 12 5 1 c
rlabel metal1 19 3 19 3 7 z
rlabel metal1 10 -19 10 -19 1 vss
rlabel polycontact -15 3 -15 3 1 a
rlabel metal1 -5 35 -5 35 5 vdd
<< end >>
