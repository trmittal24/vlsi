*nmos characteristics

.include /home/tarun/ngspice/t14y_tsmc_025_level3.txt

m1 vdd in 0 vb cmosn l=1u w=0.5u

v_dd vdd 0 3.3
v_in in 0 3.3
v_b vb 0 0

.dc v_dd 0 3.3 0.1 v_in 0 3.3 1
.dc v_in 0 3.3 0.1 v_dd 0 3.3 1


*calculating for diff width
.control

foreach iter  -2 -1 0 1
alter v_b = $iter
run
end 
.endc

*plotting diff
.control
foreach count 1 2 3 4 5 6 7 8
setplot dc$count
plot -v_dd#branch
end 
.endc

.end