* SPICE3 file created from dff.ext - technology: scmos
.include t14y_tsmc_025_level3.txt

M1000 vdd c cn vdd pfet w=9u l=2u
+ ad=348p pd=156u as=62p ps=34u 
M1001 da cn d vdd pfet w=17u l=2u
+ ad=168p pd=86u as=93p ps=52u 
M1002 vdd da d1 vdd pfet w=9u l=2u
+ ad=0p pd=0u as=133p ps=80u 
M1003 z d1 vdd vdd pfet w=9u l=2u
+ ad=117p pd=44u as=0p ps=0u 
M1004 da c z vdd pfet w=9u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1005 vdd cn cn1 vdd pfet w=9u l=2u
+ ad=0p pd=0u as=62p ps=34u 
M1006 vss c cn Gnd nfet w=5u l=2u
+ ad=228p pd=136u as=40p ps=28u 
M1007 da c d Gnd nfet w=13u l=2u
+ ad=115p pd=70u as=69p ps=44u 
M1008 da1 cn1 d1 vdd pfet w=17u l=2u
+ ad=168p pd=86u as=0p ps=0u 
M1009 vdd da1 zu vdd pfet w=9u l=2u
+ ad=0p pd=0u as=40p ps=28u 
M1010 z1 zu vdd vdd pfet w=9u l=2u
+ ad=117p pd=44u as=0p ps=0u 
M1011 da1 cn z1 vdd pfet w=9u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1012 vss da d1 Gnd nfet w=5u l=2u
+ ad=0p pd=0u as=185p ps=98u 
M1013 z d1 vss Gnd nfet w=5u l=2u
+ ad=69p pd=38u as=0p ps=0u 
M1014 da cn z Gnd nfet w=5u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1015 vss cn cn1 Gnd nfet w=5u l=2u
+ ad=0p pd=0u as=40p ps=28u 
M1016 da1 cn d1 Gnd nfet w=13u l=2u
+ ad=115p pd=70u as=0p ps=0u 
M1017 vss da1 zu Gnd nfet w=5u l=2u
+ ad=0p pd=0u as=116p ps=54u 
M1018 z1 zu vss Gnd nfet w=5u l=2u
+ ad=69p pd=38u as=0p ps=0u 
M1019 da1 cn1 z1 Gnd nfet w=5u l=2u
+ ad=0p pd=0u as=0p ps=0u 
C0 d1 vdd 11.3fF
C1 vdd da 7.1fF
C2 vss cn 3.0fF
C3 cn1 vdd 8.4fF
C4 vdd c 23.3fF
C5 cn1 vss 3.0fF
C6 zu vdd 10.4fF
C7 d1 da 2.1fF
C8 da1 vdd 7.1fF
C9 vdd cn 31.7fF
C10 z1 0 2.3fF
C11 zu 0 5.7fF
C12 vss 0 32.0fF
C13 da1 0 11.8fF
C14 cn1 0 23.9fF
C15 z 0 2.3fF
C16 d1 0 9.4fF
C17 da 0 11.6fF
C18 cn 0 45.5fF
C19 c 0 15.4fF

vdd vdd 0 5
vss vss 0 0 
v_gg_c d 0 PULSE(0 5 13n 0.1n 0.1n 25n 70n)
v_gg_d c 0 PULSE(5 0 0n 0.1n 0.1n 50n 100n)


.control
 tran 0.01n 300n
 plot (c + 10) (d + 5) zu

 .endc

.end0