*	CMOS INVERTER

.include /home/barun/vlsi/t14y_tsmc_025_level3.txt

M1 V_DS V_GS 0 0 CMOSN L = 1u W = 1u
M2 V_DS V_GS V_DD V_DD CMOSP L = 0.147u W = 1u

VDD V_DD 0 5
VIN V_GS 0 5

//VIN V_GS 0 DC 1 PULSE(0 5 1ns 0.1ns 0.1ns 2ns 4ns )
//.TRAN 0.01ns 4ns
.DC VIN 0 5 0.1 

.CONTROL
RUN
.ENDC

.CONTROL
LET V11 = DERIV(V_DS)
MEAS DC VMAX MAX V(V_DS) FROM=0ns   TO=2ns
MEAS DC VIL FIND V(V_GS) WHEN V11 = -1 FALL=LAST
PRINT 'VIL'
.ENDC

.CONTROL
FOREACH T 1 
SETPLOT DC$T
PLOT V(V_DS) V(V_GS) DERIV(V_DS)
END

.ENDC

.END
