magic
tech scmos
timestamp 1522409358
<< nwell >>
rect -2 37 80 61
<< polysilicon >>
rect 7 52 9 55
rect 19 52 21 56
rect 39 52 41 56
rect 59 52 61 56
rect 7 37 9 45
rect 7 17 9 33
rect 19 32 21 45
rect 19 17 21 28
rect 39 26 41 45
rect 59 32 61 45
rect 39 17 41 22
rect 59 17 61 28
rect 7 9 9 13
rect 19 9 21 13
rect 39 9 41 13
rect 59 9 61 13
<< ndiffusion >>
rect 3 14 7 17
rect 0 13 7 14
rect 9 13 11 17
rect 15 13 19 17
rect 21 13 39 17
rect 41 13 59 17
rect 61 13 66 17
<< pdiffusion >>
rect 0 48 7 52
rect 3 45 7 48
rect 9 48 11 52
rect 15 48 19 52
rect 9 45 19 48
rect 21 49 39 52
rect 21 45 27 49
rect 31 45 39 49
rect 41 48 48 52
rect 52 48 59 52
rect 41 45 59 48
rect 61 49 70 52
rect 61 45 66 49
<< metal1 >>
rect 11 57 70 61
rect 11 52 14 57
rect 48 52 52 57
rect -1 18 2 44
rect 8 39 13 40
rect 27 39 31 45
rect 66 39 70 45
rect 8 37 70 39
rect 11 36 70 37
rect 11 35 13 36
rect 67 17 70 36
rect 11 5 15 13
rect 11 1 71 5
<< ntransistor >>
rect 7 13 9 17
rect 19 13 21 17
rect 39 13 41 17
rect 59 13 61 17
<< ptransistor >>
rect 7 45 9 52
rect 19 45 21 52
rect 39 45 41 52
rect 59 45 61 52
<< polycontact >>
rect 7 33 11 37
rect 18 28 22 32
rect 58 28 62 32
rect 38 22 42 26
<< ndcontact >>
rect -1 14 3 18
rect 11 13 15 17
rect 66 13 70 17
<< pdcontact >>
rect -1 44 3 48
rect 11 48 15 52
rect 27 45 31 49
rect 48 48 52 52
rect 66 45 70 49
<< labels >>
rlabel metal1 35 59 35 59 5 vdd
rlabel polycontact 20 30 20 30 1 a
rlabel polycontact 60 30 60 30 1 c
rlabel metal1 40 3 40 3 1 vss
rlabel polycontact 40 24 40 24 1 b
rlabel metal1 68 34 68 34 1 zn
rlabel metal1 0 29 0 29 3 z
<< end >>
