magic
tech scmos
timestamp 1522147712
<< nwell >>
rect -28 8 60 38
<< polysilicon >>
rect -19 36 48 38
rect -19 33 -17 36
rect -5 30 -3 32
rect 17 30 19 33
rect -19 20 -17 24
rect -19 3 -17 16
rect 31 30 33 33
rect 46 30 48 36
rect -5 12 -3 13
rect -5 6 6 8
rect -19 1 -3 3
rect -19 -9 -17 1
rect -5 -1 -3 1
rect -19 -17 -17 -14
rect -5 -17 -3 -14
rect 4 -20 6 6
rect 17 -3 19 21
rect 31 14 33 21
rect 46 16 48 21
rect 32 10 33 14
rect 17 -9 19 -7
rect 31 -9 33 10
rect 46 -9 48 -3
rect 17 -16 19 -14
rect 31 -16 33 -14
rect 46 -20 48 -14
rect 4 -22 48 -20
<< ndiffusion >>
rect -10 -5 -5 -1
rect -14 -6 -5 -5
rect -23 -12 -19 -9
rect -25 -14 -19 -12
rect -17 -11 -11 -9
rect -17 -14 -16 -11
rect -12 -14 -11 -11
rect -8 -14 -5 -6
rect -3 -3 -1 -1
rect -3 -14 2 -3
rect 7 -1 8 0
rect 12 -1 13 0
rect 7 -9 13 -1
rect 7 -14 17 -9
rect 19 -14 31 -9
rect 33 -12 36 -9
rect 40 -12 46 -9
rect 33 -14 46 -12
rect 48 -12 52 -9
rect 48 -14 54 -12
rect 23 -15 27 -14
<< pdiffusion >>
rect -25 28 -19 33
rect -23 24 -19 28
rect -17 31 -16 33
rect -12 31 -11 33
rect -17 24 -11 31
rect -8 20 -5 30
rect -14 17 -5 20
rect -10 13 -5 17
rect -3 19 2 30
rect 13 28 17 30
rect 16 24 17 28
rect 13 21 17 24
rect 19 27 23 30
rect 27 27 31 30
rect 19 21 31 27
rect 33 25 46 30
rect 33 21 36 25
rect 40 21 46 25
rect 48 25 55 30
rect 48 21 53 25
rect -3 15 1 19
rect -3 13 2 15
<< metal1 >>
rect -28 35 55 38
rect 10 34 14 35
rect 23 31 26 35
rect 59 35 60 38
rect -23 25 -2 28
rect -27 -8 -24 24
rect -13 -1 -10 13
rect -5 12 -2 25
rect 8 24 12 28
rect 2 2 5 15
rect 0 1 5 2
rect -10 -5 -4 -2
rect 3 -1 5 1
rect 8 13 11 24
rect 8 10 28 13
rect 8 3 11 10
rect -7 -9 -4 -5
rect 15 -9 18 -7
rect -7 -12 18 -9
rect 36 -8 39 21
rect 53 -8 56 21
rect -16 -17 -12 -15
rect -28 -19 23 -17
rect 27 -19 60 -17
rect -28 -22 60 -19
<< ntransistor >>
rect -19 -14 -17 -9
rect -5 -14 -3 -1
rect 17 -14 19 -9
rect 31 -14 33 -9
rect 46 -14 48 -9
<< ptransistor >>
rect -19 24 -17 33
rect -5 13 -3 30
rect 17 21 19 30
rect 31 21 33 30
rect 46 21 48 30
<< polycontact >>
rect -21 16 -17 20
rect -5 8 -1 12
rect 28 10 32 14
rect 15 -7 19 -3
<< ndcontact >>
rect -27 -12 -23 -8
rect -14 -5 -10 -1
rect -16 -15 -12 -11
rect -1 -3 3 1
rect 8 -1 12 3
rect 36 -12 40 -8
rect 52 -12 56 -8
rect 23 -19 27 -15
<< pdcontact >>
rect -27 24 -23 28
rect -16 31 -12 35
rect -14 13 -10 17
rect 12 24 16 28
rect 23 27 27 31
rect 36 21 40 25
rect 53 21 57 25
rect 1 15 5 19
<< nsubstratencontact >>
rect 55 34 59 38
<< labels >>
rlabel polycontact -19 18 -19 18 1 c
rlabel metal1 -25 6 -25 6 3 cn
rlabel metal1 -12 5 -12 5 1 d
rlabel metal1 54 36 54 36 5 vdd
rlabel metal1 58 -21 58 -21 8 vss
rlabel metal1 37 4 37 4 1 z
<< end >>
